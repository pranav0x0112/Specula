package LSU;

  interface IfcLSU;
    method Action dummy();
  endinterface

  module mkLSU(IfcLSU);
    method Action dummy();
    endmethod
  endmodule

endpackage