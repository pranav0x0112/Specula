package ALU;

  interface IfcALU;
    method Action dummy();
  endinterface

  module mkALU(IfcALU);
    method Action dummy();
    endmethod
  endmodule

endpackage